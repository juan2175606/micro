magic
tech sky130A
timestamp 1652810257
<< pwell >>
rect -91 -104 20 -25
rect -90 -106 -55 -104
rect -52 -106 20 -104
<< nbase >>
rect -264 41 180 225
rect -264 40 -114 41
rect -264 39 -177 40
rect 89 39 180 41
<< nmos >>
rect -50 -98 -35 -33
<< pmos >>
rect -50 60 -35 160
<< ndiff >>
rect -90 -38 -50 -33
rect -90 -55 -81 -38
rect -64 -55 -50 -38
rect -90 -73 -50 -55
rect -90 -90 -81 -73
rect -64 -90 -50 -73
rect -90 -98 -50 -90
rect -35 -37 10 -33
rect -35 -54 -15 -37
rect 2 -54 10 -37
rect -35 -73 10 -54
rect -35 -90 -15 -73
rect 2 -90 10 -73
rect -35 -98 10 -90
<< pdiff >>
rect -95 154 -50 160
rect -95 137 -84 154
rect -67 137 -50 154
rect -95 120 -50 137
rect -95 103 -84 120
rect -67 103 -50 120
rect -95 85 -50 103
rect -95 68 -85 85
rect -68 68 -50 85
rect -95 60 -50 68
rect -35 152 9 160
rect -35 135 -15 152
rect 2 135 9 152
rect -35 116 9 135
rect -35 99 -15 116
rect 2 99 9 116
rect -35 82 9 99
rect -35 65 -15 82
rect 2 65 9 82
rect -35 60 9 65
<< ndiffc >>
rect -81 -55 -64 -38
rect -81 -90 -64 -73
rect -15 -54 2 -37
rect -15 -90 2 -73
<< pdiffc >>
rect -84 137 -67 154
rect -84 103 -67 120
rect -85 68 -68 85
rect -15 135 2 152
rect -15 99 2 116
rect -15 65 2 82
<< poly >>
rect -50 160 -35 185
rect -50 21 -35 60
rect -85 12 -35 21
rect -85 -5 -76 12
rect -59 -5 -35 12
rect -85 -13 -35 -5
rect -50 -33 -35 -13
rect -50 -123 -35 -98
<< polycont >>
rect -76 -5 -59 12
<< locali >>
rect -125 190 -64 215
rect -36 214 39 215
rect -36 190 13 214
rect -95 154 -60 190
rect -95 137 -84 154
rect -67 137 -60 154
rect -95 120 -60 137
rect -95 103 -84 120
rect -67 103 -60 120
rect -95 85 -60 103
rect -95 68 -85 85
rect -68 68 -60 85
rect -95 60 -60 68
rect -26 152 9 160
rect -26 135 -15 152
rect 2 135 9 152
rect -26 116 9 135
rect -26 99 -15 116
rect 2 99 9 116
rect -26 82 9 99
rect -26 65 -15 82
rect 2 80 9 82
rect 2 65 10 80
rect -26 60 10 65
rect -85 12 -50 21
rect -85 -5 -76 12
rect -59 -5 -50 12
rect -85 -13 -50 -5
rect -90 -38 -55 -33
rect -90 -55 -81 -38
rect -64 -55 -55 -38
rect -90 -73 -55 -55
rect -90 -90 -81 -73
rect -64 -90 -55 -73
rect -90 -128 -55 -90
rect -25 -37 10 60
rect -25 -54 -15 -37
rect 2 -54 10 -37
rect -25 -73 10 -54
rect -25 -90 -15 -73
rect 2 -90 10 -73
rect -25 -98 10 -90
rect -155 -129 13 -128
rect -127 -154 -67 -129
rect -39 -153 13 -129
rect -39 -154 40 -153
<< viali >>
rect -153 190 -125 215
rect -64 190 -36 215
rect 13 189 41 214
rect -155 -154 -127 -129
rect -67 -154 -39 -129
rect 13 -153 41 -128
<< metal1 >>
rect -166 215 50 230
rect -166 190 -153 215
rect -125 190 -64 215
rect -36 214 50 215
rect -36 190 13 214
rect -166 189 13 190
rect 41 189 50 214
rect -166 180 50 189
rect -166 -128 50 -117
rect -166 -129 13 -128
rect -166 -154 -155 -129
rect -127 -154 -67 -129
rect -39 -153 13 -129
rect 41 -153 50 -128
rect -39 -154 50 -153
rect -166 -166 50 -154
<< labels >>
rlabel metal1 -98 -142 -98 -142 1 GND
rlabel polycont -68 3 -68 3 1 A
rlabel locali -10 5 -10 5 1 Z
rlabel metal1 -84 205 -84 205 1 VDD
<< end >>
